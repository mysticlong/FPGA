//`include "src/library/DffSync_n_m.sv"
module K#(parameter n=32,m=64)(rst_i,clk_i,data_o);
input logic rst_i,clk_i;
output logic[n-1:0] data_o;
logic[n-1:0] K_i[0:m-1],K_o[0:m-1],K_shift[0:m-1];
assign           K_i[0] = 32'h428a2f98;
assign           K_i[1] = 32'h71374491;
assign           K_i[2] = 32'hb5c0fbcf;
assign           K_i[3] = 32'he9b5dba5;
assign           K_i[4] = 32'h3956c25b;
assign           K_i[5] = 32'h59f111f1;
assign           K_i[6] = 32'h923f82a4;
assign           K_i[7] = 32'hab1c5ed5;
assign           K_i[8] = 32'hd807aa98;
assign           K_i[9] = 32'h12835b01;
assign           K_i[10] = 32'h243185be;
assign           K_i[11] = 32'h550c7dc3;
assign           K_i[12] = 32'h72be5d74;
assign           K_i[13] = 32'h80deb1fe;
assign           K_i[14] = 32'h9bdc06a7;
assign           K_i[15] = 32'hc19bf174;
assign           K_i[16] = 32'he49b69c1;
assign           K_i[17] = 32'hefbe4786;
assign           K_i[18] = 32'h0fc19dc6;
assign           K_i[19] = 32'h240ca1cc;
assign           K_i[20] = 32'h2de92c6f;
assign           K_i[21] = 32'h4a7484aa;
assign           K_i[22] = 32'h5cb0a9dc;
assign           K_i[23] = 32'h76f988da;
assign          K_i[24] = 32'h983e5152;
assign          K_i[25] = 32'ha831c66d;
assign          K_i[26] = 32'hb00327c8;
assign           K_i[27] = 32'hbf597fc7;
assign           K_i[28] = 32'hc6e00bf3;
assign           K_i[29] = 32'hd5a79147;
assign           K_i[30] = 32'h06ca6351;
assign           K_i[31] = 32'h14292967;
assign           K_i[32] = 32'h27b70a85;
assign           K_i[33] = 32'h2e1b2138;
assign         K_i[34] = 32'h4d2c6dfc;
assign         K_i[35] = 32'h53380d13;
assign         K_i[36] = 32'h650a7354;
assign         K_i[37] = 32'h766a0abb;
assign         K_i[38] = 32'h81c2c92e;
assign         K_i[39] = 32'h92722c85;
assign         K_i[40] = 32'ha2bfe8a1;
assign         K_i[41] = 32'ha81a664b;
assign         K_i[42] = 32'hc24b8b70;
assign         K_i[43] = 32'hc76c51a3;
assign         K_i[44] = 32'hd192e819;
assign         K_i[45] = 32'hd6990624;
assign         K_i[46] = 32'hf40e3585;
assign         K_i[47] = 32'h106aa070;
assign         K_i[48] = 32'h19a4c116;
assign         K_i[49] = 32'h1e376c08;
assign         K_i[50] = 32'h2748774c;
assign         K_i[51] = 32'h34b0bcb5;
assign         K_i[52] = 32'h391c0cb3;
assign         K_i[53] = 32'h4ed8aa4a;
assign         K_i[54] = 32'h5b9cca4f;
assign         K_i[55] = 32'h682e6ff3;
assign         K_i[56] = 32'h748f82ee;
assign         K_i[57] = 32'h78a5636f;
assign         K_i[58] = 32'h84c87814;
assign         K_i[59] = 32'h8cc70208;
assign         K_i[60] = 32'h90befffa;
assign         K_i[61] = 32'ha4506ceb;
assign         K_i[62] = 32'hbef9a3f7;
assign         K_i[63] = 32'hc67178f2;
//dong bo
	assign K_shift[0:m-2]=K_o[1:m-1],K_shift[m-1]=K_o[0];
	DffSync_n_m#(n,m) Data_o(K_i,K_shift,rst_i,clk_i,K_o);
	assign data_o=K_o[0];
endmodule:K
 	
