module log2_x_16bit(data_i,rst_i,clk_i,Ynguyen_o,Ythapphan_o);
input logic data_i[0:15];
input logic rst_i,clk_i;
output logic[15:0] Ynguyen_o,Ythapphan_o;

logic data_io[0:15];
endmodule: log2_x_16bit

