`include "src/library/mux2to1_n.sv"
module dff_n_val#(parameter b=4,[b-1:0]val='1)(data_i,rst_i,clk_i,data_o);
	input logic [b-1:0]data_i;
	input logic	rst_i,clk_i;
	output logic[b-1:0]	data_o;
	logic[b-1:0]	data_next;
	always_ff@(posedge clk_i or negedge rst_i) begin
		if(!rst_i) data_o<=val;
		else data_o<=data_next;
	end
 mux2to1_n#(b) Q_i(data_o,data_i,rst_i,data_next);
endmodule:dff_n_val
