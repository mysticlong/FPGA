module buffer_n_m#(parameter n=32,m=64) (data_i,rst_i,clk_wr_i,clk_rd_i,data_o,fl_full)
